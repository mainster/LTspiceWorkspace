.SUBCKT 2N7292 3 2 11 V1V; REV. 6/14/90
*              D G S 
*
R21 2 1 1E9
R91 9 1 0.00654
C21 2 1 4800P
C23 2 3 200P
C24 2 4 9400P
BFDSCHRG 4 2 I=1.0*I(BVMEAS)
MOS1 4 2 1 1 MOSMOD L=1U W=1U
JFET 3 9 4 JMOD 1
DBODY 9 3 DMOD2
RSOURCE 1 10 0.01827
LSOURCE 10 11 7.5N
E41 5 11 4 1 1.0
D1 5 6 DMOD
BVPINCH 6 8 V=8.0*V(V1V)
BVMEAS 8 11 V=0*V(V1V)
DBREAK 3 7 DMOD3
BVBREAK 7 1 V=240*V(V1V)
.MODEL MOSMOD NMOS VTO=4.463 KP=12.162 TOX=1.0E+06U
.MODEL JMOD NJF VTO=-8.0 BETA=1216.2 IS=8.7E-19 RD=0.05983
.MODEL DMOD D IS=1.0E-13 N=0.03 RS=0.001
.MODEL DMOD2 D CJO=4200P TT=1000N IS=8.7E-13
.MODEL DMOD3 D IS=1.0E-13 RS=1.111 N=1.0
.ENDS