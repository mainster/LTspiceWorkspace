OP_COMP.CIR - OPAMP COMPARATOR WITH HYSTERESIS
*
VIN    1	0	SIN(0V 10VPEAK 60HZ)	
VNOISE 2	1	SIN(0V 0VPEAK 2.5KHZ)
*
* COMPARATOR
R1	2	3	1K
*R2	3	6	5K
XOP2	3 4     5	OPAMP1
RLIM	5	6	1000
D1	7	6	DZ1
D2	7	0	DZ2
*
* VREF
VREF	4	0	0V
*
*
* OPAMP MACRO MODEL, SINGLE-POLE WITH 15V OUTPUT CLAMP
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1		  1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN=100K AND POLE1=100HZ
* UNITY GAIN = DCGAIN X POLE1 = 10MHZ
EGAIN	3 0	1 2	100K
RP1	3	4	100K
CP1	4	0	0.0159UF
* ZENER LIMITER 
D1	4	7	DZ0
D2	0	7	DZ0
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
*
* 15V ZENER DIODE MODEL
.model	DZ0	D(Is=0.05u Rs=0.1 Bv=15 Ibv=0.05u)
.ENDS
*
*
* ZENER DIODE MODEL
.model	DZ1	D(Is=0.05u Rs=0.1 Bv=4.3 Ibv=0.05u)
.model	DZ2	D(Is=0.05u Rs=0.1 Bv=4.3 Ibv=0.05u)
*
* ANALYSIS
.TRAN 	0.1MS 34MS
*
* VIEW RESULTS
.PRINT TRAN	V(2) V(6)
.PROBE
.END