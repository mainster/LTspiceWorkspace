*==========================================================
* Analog Devices Linear ICs
*
* This model was developed by:
* AEI Systems, LLC
* 5777 W. Century Blvd. Suite 876
* Los Angeles, California 90045
* Copyright 2002, all rights reserved.
*
* This model is subject to change without notice.
* Users may not directly or indirectly re-sell or 
* re-distribute this model.
*
* For more information contact 
* AEi by email: info@aeng.com. http://www.AENG.com
*
*==========================================================
***************
* |=======================================================
* | ADI VARIABLE GAIN AMPLIFIER MACRO-MODEL AD8331/2/4 LNA
* |=======================================================
*
* Connections:
*
.SUBCKT VGA VIP VIN MODE GAIN VCM RCLMP HILO VPOS VOH VOL COMM ENBV
EB2 35 0 Value = {10**(V(GAIN1)*2.5-2.5)}
R36 POST1 0 1MEG
GB7 59 0 Value = {I(VSNS4)*V(ENV1)}
GB8 52 0 Value = {I(VSNS3)*V(ENV1)}
GB3 0 39 Value = {(V(VIP)-V(VIN))*V(GAIN2)*10U}
R27 VIP MID1 100
R28 VIN MID1 100
R29 GAIN COMM 10MEG
R19 VOL COMM 1MEG
R33 39 0 1MEG
EB1 37 0 Value = {IF(V(MODE) - V(COMM) < 1.625 , V(GAIN) - V(COMM) , 1.04 - V(GAIN) + V(COMM))}
E4 MID1 COMM VPOS COMM 0.5
R30 MODE COMM 200K
R31 37 GAIN1 1K
C4 GAIN1 0 217P
R10 VCM MID1 30
R37 HILO COMM 50K
EB4 HILO1 0 Value = {V(HILO2) * (5.9566 - 1.4962) + 1.4962}
R38 48 HILO2 1K
C5 HILO2 0 10P
GB5 0 POST1 Value = {V(VGA1)*V(HILO1)*V(ENV1)*0.1U}
G2 MID1 68 0 POST1 0.5U
R52 68 MID1 1MEG
EB14 48 0 Value = {IF(V(HILO) - V(COMM) < 1.625 , 0 , 1)}
EB15 CLMP1 0 Value = {V(CLMP2) - 0.36 + 0.12*V(HILO2) - 0.12}
D29 36 GAIN2 _DLIM2 
VSNS4 71 72 DC=0
R56 72 VOL 1
F7 VPOS 71 VLP4 -1
F8 71 COMM VLN4 -1
VLN4 0 60 DC=.63
D20 57 59 _DDEF 
D22 59 62 _DDEF 
D21 59 61 _DDEF 
D19 56 59 _DDEF 
R50 58 57 100
R51 60 61 100
VLP4 58 0 DC=.63
V14 62 0 DC=4.36
R54 VPOS VOL 100MEG
R55 VOL COMM 100MEG
R53 68 71 100MEG
V13 0 56 DC=4.36
E8 MID1 69 CLMP1 0 0.25
D26 69 68 _DLIM 
D25 68 70 _DLIM 
E9 70 MID1 CLMP1 0 0.25
I6 COMM VPOS DC=236.1U
G1 MID1 64 POST1 0 0.5U
R45 64 MID1 1MEG
VSNS3 66 67 DC=0
R49 67 VOH 1
F5 VPOS 66 VLP3 -1
F6 66 COMM VLN3 -1
VLN3 0 53 DC=.63
D16 50 52 _DDEF 
D18 52 55 _DDEF 
D17 52 54 _DDEF 
D15 49 52 _DDEF 
R43 51 50 100
R44 53 54 100
VLP3 51 0 DC=.63
V12 55 0 DC=4.36
R47 VPOS VOH 100MEG
R48 VOH COMM 100MEG
R46 64 66 100MEG
V11 0 49 DC=4.36
E10 MID1 63 CLMP1 0 0.25
D24 63 64 _DLIM 
D23 64 65 _DLIM 
E11 65 MID1 CLMP1 0 0.25
R57 RCLMP COMM 10.7235K
C3 VGA1 0 1.061F
R34 VGA1 42 1MEG
D27 40 39 _DLIM 
I7 COMM RCLMP DC=233.13U
E14 CLMP2 0 73 0 2
V15 0 40 DC=5
E13 73 0 RCLMP COMM 0.98625
R41 ENBV COMM 70K
EB6 75 0 Value = {IF(V(ENBV) - V(COMM) < 1.625 , 0 , 1)}
R42 75 ENV1 1K
C7 ENV1 0 10P
R18 VOH COMM 1MEG
G3 VPOS COMM ENV1 0 14M
D28 39 41 _DLIM 
V16 41 0 DC=5
E5 42 0 39 0 11.22
R35 43 44 1MEG
VSR1 42 43 DC=0
F9 VGA1 0 VSR1 1
E12 47 0 VGA1 0 1
D31 44 46 _DLIM 
V19 46 47 DC=2.01
D32 45 44 _DLIM 
V20 47 45 DC=2.01
V17 36 0 DC=0.004
D30 GAIN2 38 _DLIM 
V18 38 0 DC=0.9
R32 GAIN2 35 1K
.MODEL _DDEF D
.MODEL _DLIM D EG=.222 N=.2
.MODEL _DLIM2 D EG=.222 N=.0002
.ENDS
