DG4
*SPICE_NET
.INCLUDE DG_MOS.LIB
.TRAN .1N 1000N 800N
.lib standard.dio
*ALIAS  V(7)=TANK
*ALIAS  V(2)=DRAIN
*ALIAS  V(5)=VG2
*ALIAS  V(8)=VG1
.PRINT TRAN  V(7)  V(2)  V(5)  V(8) 
.PRINT TRAN  V(10) 
R1 1 4 270
R2 3 2 100
C1 1 4 .05U
C2 2 0 .05U
R3 3 5 180K
V1 3 0 18
R4 5 10 20K
R5 5 5 50K
R6 5 0 50K
R7 8 0 47K
D1 8 0 1N914
C3 7 0 10P
L1 7 4 .2024U
L2 4 0 .0506U
C4 7 8 47P
C5 5 0 .01U
V2 10 0 PULSE 0 7 0 0 0 50N 100N
X1 2 5 8 1 MN201 
.END
