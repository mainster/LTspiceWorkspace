* D:\LTspiceWorldTour2009\SubcktMOSFET.asc
V1 N001 0 0
V2 N002 0 0
XM2 N001 N002 0 IRF_7401
.dc V1 0 20 10m V2 2 14 2
.SUBCKT IRF_7401 1 2 3
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 Is=1e-32 Vto=1.3 Lambda=.0087315 KP=124 Cgso=1.4e-5 Cgdo=1.4e-06
RS 8 3 0.0153334
D1 3 1 MD
.MODEL MD D Is=10n Rs=63m N=1.36 BV=20 IBV=250u EG=1 XTI=3 TT=100n Cjo=1n Vj=5 M=.72 FC=.5
RDS 3 1 16Meg
RD 9 1 1.9m
RG 2 7 9.481
D2 4 5 MD1
.MODEL MD1 D Is=1e-32 N=50 Cjo=2.15n Vj=.526 M=0.744 Fc=1e-8
D3 0 5 MD2
.MODEL MD2 D Is=1e-10 N=.4 Rs=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3n
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
.MODEL MD3 D Is=1e-10 N=.4
.ENDS IRF_7401
.backanno
.end
