DGYFS
.OPTIONS LIMPTS=2000 ITL2=100
*OPT VTEMP=0 TO 3 STEP=1
*OPT TEMP=-.5 TO 1.5 STEP=.2
*.AC DEC 10 1K 10K
.DC VDS 0 10 .1 VGS1 -1.5 1 .5
************
*SPICE_NET
.INCLUDE DG_MOS.LIB
*ALIAS  I(V2)=ID
*ALIAS  V(1)=YFS
.PRINT AC I(V2) IP(V2) V(1)  VP(1) V(4)
.PRINT DC I(V2)
VDS 2 0 15
RDS 1 5 1
VGS2 3 0 4
*VTEMP
VGS1 4 0 
*TEMP AC 1
R2 4 0 1MEG
V2 2 5 
X1 1 3 4 0 MN201
.END
