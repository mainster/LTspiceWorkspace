DG3
*SPICE_NET
.INCLUDE DG_MOS.LIB
.TRAN .05N 20N
*.AC DEC 10 100K 1000MEG
*ALIAS  V(11)=OUTPUT
*ALIAS  V(1)=INPUT
*ALIAS  V(2)=VIN
.PRINT AC  V(11)  VP(11)  V(1)  VP(1) 
.PRINT AC  V(2)  VP(2) 
.PRINT TRAN  V(11)  V(1)  V(2) 
L1 2 3 1M
C1 12 2 5P
C2 3 0 500P
R1 0 3 300K
R2 3 7 360K
R3 7 6 820K
C3 6 0 500PF
L2 6 9 1M
C4 2 0 4P
X1 9 7 2 8 MN201 
C5 7 0 500P
R5 8 0 270
C6 8 0 500P
C7 9 0 5P
R6 11 0 50
C8 9 11 5P
R7 1 12 50
V2 6 0 8
V1 1 0 SIN 0 10 200MEG AC 1
.END
