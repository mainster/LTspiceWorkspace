* C:\data\Ltc_Spice\Infineon SPD22N08S2L\infineon_xnmos5_test.asc
R1 N002 N001 10
XU1 out N001 0 N004 N005 SPD22N08S2L-50
V1 N003 0 10
R2 N003 out 10
V2 N002 0 PULSE(0 5 10n 5n 5n 200n 1000n)
R3 N005 0 1
.tran 0 4u 0 5n
.INCLUDE SPD22N08S2L.sub
.PROBE  
* .include optimos_n.lib
* Watch V(out)!
.end
