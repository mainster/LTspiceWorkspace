* D:\Arrow\2N5817.asc
V1 0 N001 0
Q1 N001 N002 0 0 2N5817
I1 N002 0 0
.dc V1 0 3 1m I1 20u 100u 20u
.model 2N5817  PNP(Is=650.6E-18 Xti=3 Eg=1.11 Vaf=115.7 Bf=127 Ne=1.829
+                               Ise=99.99f Ikf=1.079 Xtb=1.5 Br=3.752 Nc=2 Isc=0 Ikr=0 Rc=.715
+                               Cjc=14.76p Mjc=.5383 Vjc=.75 Fc=.5 Cje=19.82p Mje=.3357 Vje=.75
.end
