Simple SC integrator

.param supply=3

vphi1   phi1   0 pulse({supply} 0  530ns 180ps 180ps 503ns 1u)
vphi1i  phi1i  0 pulse(0 {supply}  530ns 180ps 180ps 503ns 1u)
vphi2   phi2   0 pulse(0 {supply}  560ns 180ps 180ps 497ns 1u)
vphi2i  phi2i  0 pulse({supply} 0  560ns 180ps 180ps 497ns 1u)

.subckt switch a avdd avss c xc z
mmp z xc a avdd p1 w=3u l=0.6u ad=40.5p as=40.5p
+pd=62.7u ps=62.7u nrd=26.67m nrs=26.67m
mmn a c z avss n1 w=1.5u l=0.6u ad=20.25p as=20.25p
+pd=32.7u ps=32.7u nrd=53.33m nrs=53.33m
.ends switch

.subckt ota avdd avss ibp vin vip vo
mm4 net9 vip sp sp p1 w=90u l=1.8u ad=121.5p as=121.5p
+pd=182.7u ps=182.7u nrd=8.889m nrs=8.889m
mm3 gn vin sp sp p1 w=90u l=1.8u ad=121.5p as=121.5p
+pd=182.7u ps=182.7u nrd=8.889m nrs=8.889m
rrc net9 net4 5k
ccc net4 vo 1.5p
mm7 vo net9 avss avss n1 w=45u l=1.5u ad=60.75p as=60.75p
+pd=92.7u ps=92.7u nrd=17.78m nrs=17.78m
mm6 net9 gn avss avss n1 w=18u l=4u ad=24.3p as=24.3p
+pd=38.7u ps=38.7u nrd=44.44m nrs=44.44m
mm5 gn gn avss avss n1 w=18u l=4u ad=24.3p as=24.3p
+pd=38.7u ps=38.7u nrd=44.44m nrs=44.44m
mm2 vo ibp avdd avdd p1 w=15u l=1u ad=20.25p as=20.25p
+pd=32.7u ps=32.7u nrd=53.33m nrs=53.33m m=10
mm1 sp ibp avdd avdd p1 w=15u l=1u ad=20.25p as=20.25p
+pd=32.7u ps=32.7u nrd=53.33m nrd=53.33m m=3
mm0 ibp ibp avdd avdd p1 w=15u l=1u ad=20.25p as=20.25p
+pd=32.7u ps=32.7u nrd=53.33m nrs=53.33m
.ends ota

vdd avdd 0 dc {supply}
vss avss 0 dc 0
vcm vcm 0 dc 1
vin vin vcm dc 0 sin(0 0.3 20k)

xs1 vin avdd avss phi1 phi1i c1n switch
c1 c1n c1p 0.2p
xs2 c1p avdd avss phi2 phi2i vin_ota switch
xs3 vcm avdd avss phi2 phi2i c1n switch
xs4 c1p avdd avss phi1 phi1i vcm switch
c2 vin_ota vo 1p
xota avdd avss ibp vin_ota vcm vo ota
ibias avdd ibp -3.9u

.model n1 nmos level=8
+ Tnom=27.0
+ nch= 1.024685E+17  tox=1.00000E-08 xj=1.00000E-07
+ lint= 3.75860E-08 wint=-2.02101528644562E-07
+ vth0= .6094574   k1= .5341038  k2= 1.703463E-03  k3=-17.24589
+ dvt0= .1767506  dvt1= .5109418  dvt2=-0.05
+ nlx= 9.979638E-08  w0=1e-6
+ k3b= 4.139039
+ vsat= 97662.05  ua=-1.748481E-09  ub= 3.178541E-18  uc=1.3623e-10 
+ rdsw= 298.873  u0= 307.2991 prwb=-2.24e-4
+ a0= .4976366
+ keta=-2.195445E-02  a1= .0332883  a2= .9
+ voff=-9.623903E-02  nFactor= .8408191  cit= 3.994609E-04
+ cdsc= 1.130797E-04
+ cdscb=2.4e-5
+ eta0= .0145072  etab=-3.870303E-03
+ dsub= .4116711
+ pclm= 1.813153  pdiblc1= 2.003703E-02  pdiblc2= .00129051 pdiblcb=-1.034e-3
+ drout= .4380235  pscbe1= 5.752058E+08  pscbe2= 7.510319E-05
+ pvag= .6370527 prt=68.7 ngate=1.e20 alpha0=1.e-7 beta0=28.4 
+ prwg=-0.001 ags=1.2
+ dvt0w=0.58 dvt1w=5.3e6 dvt2w=-0.0032
+ kt1=-.3  kt2=-.03
+ at= 33000
+ ute=-1.5
+ ua1= 4.31E-09  ub1= 7.61E-18  uc1=-2.378e-10
+ kt1l=1e-8
+ wr=1 b0=1e-7 b1=1e-7 dwg=5e-8 dwb=2e-8 delta=0.015
+ cgdl=1e-10 cgsl=1e-10 cgbo=1e-10 xpart=0.0
+ cgdo=0.4e-9 cgso=0.4e-9 
+ clc=0.1e-6
+ cle=0.6
+ ckappa=0.6

.model p1 pmos level=8
+ Tnom=27.0
+ nch= 5.73068E+16  tox=1.00000E-08 xj=1.00000E-07
+ lint= 8.195860E-08 wint=-1.821562E-07
+ vth0= -.86094574   k1= .341038  k2= 2.703463E-02  k3=12.24589
+ dvt0= .767506  dvt1= .65109418  dvt2=-0.145
+ nlx= 1.979638E-07  w0=1.1e-6
+ k3b= -2.4139039
+ vsat= 60362.05  ua=1.348481E-09  ub= 3.178541E-19  uc=1.1623e-10 
+ rdsw= 498.873  u0= 137.2991 prwb=-1.2e-5
+ a0= .3276366
+ keta=-1.8195445E-02  a1= .0232883  a2= .9
+ voff=-6.623903E-02  nFactor= 1.0408191  cit= 4.994609E-04
+ cdsc= 1.030797E-3
+ cdscb=2.84e-4
+ eta0= .0245072  etab=-1.570303E-03
+ dsub= .24116711
+ pclm= 2.6813153  pdiblc1= 4.003703E-02  pdiblc2= .00329051 pdiblcb=-2.e-4
+ drout= .1380235  pscbe1= 0  pscbe2=1.e-28 
+ pvag= -.16370527
+ prwg=-0.001 ags=1.2
+ dvt0w=0.58 dvt1w=5.3e6 dvt2w=-0.0032
+ kt1=-.3  kt2=-.03 prt=76.4
+ at= 33000
+ ute=-1.5
+ ua1= 4.31E-09  ub1= 7.61E-18  uc1=-2.378e-10
+ kt1l=0
+ wr=1 b0=1e-7 b1=1e-7 dwg=5e-8 dwb=2e-8 delta=0.015
+ cgdl=1e-10 cgsl=1e-10 cgbo=1e-10 xpart=0.0
+ cgdo=0.4e-9 cgso=0.4e-9 
+ clc=0.1e-6
+ cle=0.6
+ ckappa=0.6
.tran 0 100u 0 1u
