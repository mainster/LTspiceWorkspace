* D:\Test_lt\BLF245_pspice.asc
L1 N009 2 24.5nh
C1 0 N003 100pF
C2 N002 0 30p
C3 N002 Vin 20p
R1 1 N003 1K
L3 N005 2 98nH
C5 0 N005 100pF
C6 N005 N008 100nF
C7 N009 Vout 18pF
C8 N009 Vout 30p
L4 N005 N006 70mh
R3 0 N008 10
C9 Vout 0 27pF
C10 Vout 0 24pF
Rload Vout 0 50
L2 1 N002 13.5nh
Rgen N001 Vin 50
V1 N001 0 SIN(0 510m 50Meg) AC 1
R6 N006 N007 1
R7 N003 N004 1
C4 0 N003 100n
V2 N004 0 0
V3 N007 0 0
.tran 0 1u 0 .1n
.include BLF245_28V_50MA.l2P
X1 1 2 0 BLF245_28V_50MA
.probe
* .ac dec 100 1e6 1e9
*.backanno
.end
