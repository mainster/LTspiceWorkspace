ADA4700 SPICE Macro-model      
* Description: Amplifier
* Generic Desc: 10V/100V, BIPOLAR
* Developed by: DB / ADSJ
* Revision History: 
*02/18/2014 - initial release
*02/26/2014 rev 0.1 - Edited subckt line
* 0.1 (02/2014)
*
* Copyright 2014 by Analog Devices
*
* T=25�C
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.

*****************************************************
*                      in+ in- vps+ vps- out
.SUBCKT ADA4700  1   2   99   50   5
*
*****************************************************
*
*****************************************************
* input gm (voltage -> current) stage
q1    99      3       6      50        npn1  10
q2    99      4       7      50        npn1  10
q3    50      3       6      50        pnp1   1
q4    50      4       7      50        pnp1   1
c3    1       50      5.0pf
c4    2       50      5.0pf
c5    3       4       0.5pf
r5    1       3       2k
r6    2       4       2k
d01   6       8       d1
d02   7       9       d1
d03   9       8       d1
d04   8       9       d1
g01   8       50      56       55     160e-6
g02   9       50      56       55     160e-6
e01   10      55      87       9      1.00
e02   91      55      11       55     1.00
e03   92      55      12       55     1.00
e04   93      91      56       55     12e-3
e05   92      94      56       55     12e-3
d05   10      11      d1
d06   12      10      d1
d07   95      93      d1
d08   94      96      d1
r7    55      95      200
r8    96      55      200
g04   55      14      55       95     3.00e-3
g05   15      55      96       55     3.00e-3
g06   11      14      56       55     100e-6
g07   15      12      56       55     100e-6
*
* input (NPN) base current caneclation
q5    99      45      44      50        npn1  10
g14   44      50      56      55        160e-6
e15   99      46      56      55        0.6
g20   99      45      46      45        10e-6
g21   99      3       46      45        10e-6
g22   99      4       46      45        10e-6
*
********************************************************
* current mirror, voltage gain, and compensation at negative supply
g08   14      50      14     50        0.5e-3
g09   18      50      14     50        0.5e-3
c13   16      20      3.0pf
c15   20      18      15pf
c17   14      50      4.0pf
c19   20      50      3.0pf
r13   14      16      2.0k
c22   18      50      6.0pf
c23   21      50      20pf
r10   14      50      1e9
r21   18      50      400e6
*
********************************************************
* current mirror, voltage gain, and compensation at postive supply
g10   99      15      99      15      0.5e-3
g11   99      19      99      15      0.5e-3
c14   17      20      3.0pf
c16   20      19      15pf
c18   99      15      4.0pf
c20   99      20      3.0pf
r14   15      17      2.0k
c24   19      99      6.0pf
c25   22      99      20pf
r11   99      15      1e9
r23   19      99      400e6
*
********************************************************
* unit gain voltage buffer and output drive and bias
q12   34      34      29      50        pnp1  600
q13   35      35      29      50        npn1  300
e06   28      50      27      50        1.0
d9    23      21      d1
d10   24      23      d1
d11   20      24      d1
d12   25      20      d1
d13   26      25      d1
d14   22      26      d1
d15   32      27      d1
d16   27      33      d1
d21   34      29      d1
d22   29      35      d1
r15   21      18      1.2k
r16   19      22      1.2k
r19   20      21      7.0k
r20   22      20      7.0k
r27   29      28      2.0k
* noiseless 40k resistors
g18   20      27      20      27      25e-6
*
g12   34      50      56      55     100e-6
g13   99      35      56      55     100e-6
e13   32      50      54      55     2.6
e14   99      33      54      55     2.7
*
* output transistors w/short current limit and output feedback compensation
q17   99      37      39      50        npn1  300
q18   50      36      38      50        pnp1  600
q19   43      39      38      50        npn1  1
q20   42      38      39      50        pnp1  1
d19   22      43      d1
d20   42      21      d1
r3    39      5       20
r4    5       38      20
r17   35      37      2.0k
r18   34      36      1.0k
* current boost for output transistors
g16   36      50      36      34      15e-3
g17   99      37      35      37      3.0e-3
*
r25   42      21      100k
r26   22      43      100k
*
c1    5       41      20.0pf
r1    22      41      5.0k
c2    5       40      20.0pf
r2    21      40      5.0k
*
********************************************************
* macromodel turn on control and bias
*
* Generate 1.0 volt reference
qb1   60      60      99      50      pnp1   1
qb2   62      61      50      50      npn1   1
qb3   64      62      63      50      npn1   10
d64   65      64      d1
d65   99      65      d1
d66   66      64      d1
d67   67      55      d1
d68   68      55      d1
rb1   60      61      2e6
rb2   61      62      1.0k
rb3   61      50      500k
rb4   63      50      300
rb5   65      64      20k
rb6   99      65      20k
rb7   99      66      20k
rb8   67      55      10e6
rb9   68      55      160e6
g67   99      67      99      66     160e-6
g68   99      68      99      66     10e-6
e67   69      55      67      55     0.77
e68   70      69      67      68     7.90
*
* Buffer and filter 1.0 volt reference
r51   70      51      10k
c51   51      55      40pf
e51   53      55      51      55     1.00
r52   53      52      10k
c52   52      55      40pf
e52   56      55      52      55     1.00
*
* Generate voltage half way between the power suppplies
eb1   55      50      99      50     0.50
*
* Generate  one diode voltage 
g54   55      54      56      55     100e-6
d40   54      55      d1
rb10  54      55      20k
*
********************************************************
* input error adjusts and input noise
*
* Vos
e84   84      8       56      55     1e-15
*
* Input Voltage Noise flat band and 1/f
e87   87      84      78      79     1.6
d76   76      55      dnoise
d77   77      55      dnoise
g76   55      76      56      55     160e-6
g77   55      77      56      55     160e-6
c77   79      78      5.0pf
r77   79      78      2.0k
r78   76      78      300k
r79   77      79      300k
*
* Input Current Noise flat band and 1/f
d80   80      55      dnoise
d81   81      55      dnoise
d82   82      55      dnoise
g80   55      80      56      55     160e-6
g81   55      81      56      55     160e-6
g82   55      82      56      55     160e-6
g31   2       50      81      80     0.20e-6
g32   1       50      82      80     0.20e-6
*
********************************************************
* adjust supply current
*
* set supply current at low voltage supply voltage
g15   99      50      56      55     600e-6
*
* set supply current change with supply voltage change
r30   99      50      1.0e6
*
********************************************************
* esd diodes
d51   50      1       d2
d52   1       99      d2
d53   50      2       d2
d54   2       99      d2
d55   50      5       d2
d56   5       99      d2
d57   50      99      dz120
*
********************************************************
* models
*
.MODEL npn1 NPN is=1e-16, bf=200, vaf=150, ikf=100e-6
*.MODEL npn1 NPN is=1e-16, bf=400, vaf=150, ikf=100e-6
.MODEL pnp1 PNP is=1e-16, bf=100, vaf=100, ikf=50e-6
*
*.model d1     d  is=1e-14, rs=1.0
.model d1     d  is=1e-14, rs=10
.model d2     d  is=1e-14, rs=1.0
.model dnoise d  is=1e-14, rs=1.0, kf=5.0e-11
.model dz120  d  is=1e-13, rs=1.0, bv=120, ibv=5e-4
*
********************************************************
* generator format
* g_gen  out_sink  out_source  input_pos  input_neg  gain(amp/volt)
* e_gen  out_pos   out_neg     input_pos  input_neg  gain(volt/volt)
********************************************************
*
.ENDS ADA4700
*
*****************************************************
