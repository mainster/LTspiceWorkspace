* Z:\home\mainster\CODES_local\LTSpice_projects\diskret_op\diskret_op_minimal.asc
Q1 Vo- in- N001 0 PNP1
Q2 Vo+ in+ N001 0 PNP1
I1 V+ N001 25u load
I2 V+ N002 200u
Q3 Vo- Vo- V- 0 NPN1
Q4 Vo+ Vo- V- 0 NPN1
XIdv N005 Vo+ arrow_curr arrow_curr Rsh=1m
Q5 V+ N003 N006 0 NPN1
Q6 N002 N006 V- 0 NPN1
I4 N006 V- 20u
Q7 V+ N002 out 0 NPN1
Q8 V- N002 out 0 PNP1
C1 N002 N003 {Ccomp}
XU1 V+ vdc_single V={VCC}
XU2 V- vdc_single V={VEE}
V1 in+ 0 SINE(0 10m 1k 5m) AC 1
R2 N005 0 100k
R1 0 0 100meg
E1 in- 0 in+ 0 -1
R3 Vo- V- 50t
.model NPN NPN
.model PNP PNP
.lib C:\Program Files (x86)\LTC_ALL\LTspiceIV_4.18_multiLibs\lib\cmp\standard.bjt
.model NPN1 npn (IS=4.679E-14 Bf=Bfn)
.model PNP1 pnp (IS=4.679E-14 Bf={BFp})
.model NPN11 npn (Is={I0/exp(0.6/26m)} Bf=400)
.model PNP11 pnp (Is={I0/exp(0.6/26m)} Bf=300)
.param I0=100u
.param Ccomp=30p
.param VCC=30V
.param VEE=-30V
* .tran 10m
.dc V1 -150m 150m 1m
* plot:\n-------\nIx(Idv:out)\n-40u/(4*26m)*V(in+,in-)/(1V/1A)*0.5*(sgn(V(in+,in-)+80m)-sgn(V(in+,in-)-80m))\nd( -40u/(4*26m)*V(in+,in-)/(1V/1A)*0.5*(sgn(V(in+,in-)+80m)-sgn(V(in+,in-)-80m)) )
* .model PNP1 PNP(IS=3.83E-14 NF=1.008 ISE=1.22E-14 NE=1.528 BF=344.4 IKF=0.08039 VAF=21.11 NR=1.005 ISC=2.85E-13 NC=1.28 BR=14.84 IKR=0.047 VAR=32.02 RB=1 IRB=1.00E-06 RBM=1 RE=0.6202 RC=0.5713 XTB=0 EG=1.11 XTI=3 CJE=1.23E-11 VJE=0.6106 MJE=0.378 TF=5.60E-10 XTF=3.414 VTF=5.23 ITF=0.1483 PTF=0 CJC=1.08E-11 VJC=0.1022 MJC=0.3563 XCJC=0.6288 TR=1.00E-32 CJS=0 VJS=0.75 MJS=0.333 FC=0.8027 Vceo=45 Icrating=100m mfg=Philips)\n.model NPN1 NPN(IS=2.39E-14 NF=1.008 ISE=3.545E-15 NE=1.541 BF=294.3 IKF=0.1357 VAF=63.2 NR=1.004 ISC=6.272E-14 NC=1.243 BR=7.946 IKR=0.1144 VAR=25.9 RB=1 IRB=1.00E-06 RBM=1 RE=0.4683 RC=0.85 XTB=0 EG=1.11 XTI=3 CJE=1.358E-11 VJE=0.65 MJE=0.3279 TF=4.391E-10 XTF=120 VTF=2.643 ITF=0.7495 PTF=0 CJC=3.728E-12 VJC=0.3997 MJC=0.2955 XCJC=0.6193 TR=1.00E-32 CJS=0 VJS=0.75 MJS=0.333 FC=0.9579 Vceo=45 Icrating=100m mfg=Philips)
.param Bfn=400
.param Bfp=300
.param alpha=Bfn/(Bfn+1)
.lib EIT_sub/vdc_single.sub
.lib MDB_sub/arrow_curr.sub
.backanno
.end
