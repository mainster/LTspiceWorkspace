BUCK_BASIC.CIR - BASIC BUCK CONVERTER
*
* SWITCH DRIVER 
VCTRL	10	0	PULSE(0V 5V 0 0.01US 0.01US 5US 20US)
R10	10	0	1MEG
*
* INPUT VOLTAGE
VIN	1	0	DC	20
*
* CONVERTER
SW1	1 2	10 0 	SW
D1	0	2	DSCH
L1	2	3	50UH
C1	3	0	25UF
*
* LOAD
RL	3	0	5
*
*
.MODEL	SW	VSWITCH(VON=5V VOFF=0V RON=0.01 ROFF=1MEG)
.MODEL DSCH D( IS=0.0002 RS=0.05 CJO=5e-10  )
*
* ANALYSIS
.TRAN 	1US  	800US
*.TRAN 	0.1US  	840US  800US 0.1US
*
* VIEW RESULTS
.PLOT	TRAN	V(2) V(3)
.PROBE
.END